force -freeze /E 0000 0 ns, 0001 20 ns, 0010 40 ns, 0011 60 ns -r 80 ns